library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity lut_core is
    Generic (
        num_rows : integer :=128;
        num_cols : integer :=128;
        num_theta_angles : integer := 216;
        num_phi_angles : integer :=3
    );
  Port ( 
    clk : in std_logic;
    requested_row : in integer;
    requested_col : in integer;
    requested_theta : in integer;
    requested_phi : in integer;
    necessary_voltage_psi0 : out integer range 0 to 255;
    necessary_voltage_psi1 : out integer range 0 to 255;
    necessary_voltage_psi2 : out integer range 0 to 255;
    necessary_voltage_psi3 : out integer range 0 to 255;
    necessary_voltage_psi4 : out integer range 0 to 255;
    returned_theta_ang : out integer
  );
end lut_core;

architecture Behavioral of lut_core is

type voltage_LUT is array (num_rows-1 downto 0, num_cols-1 downto 0, num_theta_angles-1 downto 0, num_phi_angles-1 downto 0) of integer range 0 to 255;
type theta_LUT is array (num_theta_angles-1 downto 0) of integer;

constant psi0_volt_LUT : voltage_LUT :=(
(15 => (7 => (0 => (others => 7), 
1 => (others => 8), 
2 => (others => 8), 
3 => (others => 9), 
4 => (others => 10), 
5 => (others => 11), 
6 => (others => 12), 
7 => (others => 13), 
8 => (others => 14), 
9 => (others => 14), 
10 => (others => 15), 
11 => (others => 16), 
12 => (others => 17), 
13 => (others => 18), 
14 => (others => 18), 
15 => (others => 19), 
16 => (others => 2), 
17 => (others => 3), 
18 => (others => 4), 
19 => (others => 4), 
20 => (others => 5), 
21 => (others => 6), 
22 => (others => 7), 
23 => (others => 7), 
24 => (others => 7), 
25 => (others => 8), 
26 => (others => 9), 
27 => (others => 10), 
28 => (others => 10), 
29 => (others => 11), 
30 => (others => 12), 
31 => (others => 12), 
32 => (others => 13), 
33 => (others => 13), 
34 => (others => 13), 
35 => (others => 16), 
36 => (others => 16), 
37 => (others => 17), 
38 => (others => 18), 
39 => (others => 19), 
40 => (others => 19), 
41 => (others => 20), 
42 => (others => 21), 
43 => (others => 22), 
44 => (others => 22), 
45 => (others => 9), 
46 => (others => 10), 
47 => (others => 11), 
48 => (others => 12), 
49 => (others => 13), 
50 => (others => 14), 
51 => (others => 15), 
52 => (others => 16), 
53 => (others => 17), 
54 => (others => 18), 
55 => (others => 19), 
56 => (others => 20), 
57 => (others => 21), 
58 => (others => 28), 
59 => (others => 29), 
60 => (others => 30), 
61 => (others => 31), 
62 => (others => 32), 
63 => (others => 33), 
64 => (others => 34), 
65 => (others => 34), 
66 => (others => 35), 
67 => (others => 36), 
68 => (others => 37), 
69 => (others => 38), 
70 => (others => 39), 
71 => (others => 40), 
72 => (others => 88), 
73 => (others => 89), 
74 => (others => 90), 
75 => (others => 91), 
76 => (others => 92), 
77 => (others => 92), 
78 => (others => 93), 
79 => (others => 105), 
80 => (others => 106), 
81 => (others => 107), 
82 => (others => 108), 
83 => (others => 109), 
84 => (others => 110), 
85 => (others => 111), 
86 => (others => 112), 
87 => (others => 113), 
88 => (others => 114), 
89 => (others => 115), 
90 => (others => 116), 
91 => (others => 116), 
92 => (others => 122), 
93 => (others => 123), 
94 => (others => 124), 
95 => (others => 125), 
96 => (others => 125), 
97 => (others => 126), 
98 => (others => 127), 
99 => (others => 128), 
100 => (others => 129), 
101 => (others => 130), 
102 => (others => 131), 
103 => (others => 131), 
104 => (others => 132), 
105 => (others => 133), 
106 => (others => 134), 
107 => (others => 119), 
108 => (others => 120), 
109 => (others => 121), 
110 => (others => 122), 
111 => (others => 123), 
112 => (others => 124), 
113 => (others => 125), 
114 => (others => 126), 
115 => (others => 115), 
116 => (others => 115), 
117 => (others => 116), 
118 => (others => 116), 
119 => (others => 117), 
120 => (others => 118), 
121 => (others => 119), 
122 => (others => 120), 
123 => (others => 121), 
124 => (others => 122), 
125 => (others => 123), 
126 => (others => 124), 
127 => (others => 124), 
128 => (others => 125), 
129 => (others => 126), 
130 => (others => 145), 
131 => (others => 146), 
132 => (others => 147), 
133 => (others => 147), 
134 => (others => 148), 
135 => (others => 149), 
136 => (others => 150), 
137 => (others => 150), 
138 => (others => 151), 
139 => (others => 152), 
140 => (others => 153), 
141 => (others => 153), 
142 => (others => 154), 
143 => (others => 155), 
144 => (others => 156), 
145 => (others => 156), 
146 => (others => 156), 
147 => (others => 158), 
148 => (others => 159), 
149 => (others => 160), 
150 => (others => 161), 
151 => (others => 176), 
152 => (others => 177), 
153 => (others => 178), 
154 => (others => 179), 
155 => (others => 180), 
156 => (others => 181), 
157 => (others => 182), 
158 => (others => 183), 
159 => (others => 184), 
160 => (others => 185), 
161 => (others => 185), 
162 => (others => 186), 
163 => (others => 187), 
164 => (others => 188), 
165 => (others => 188), 
166 => (others => 186), 
167 => (others => 187), 
168 => (others => 188), 
169 => (others => 236), 
170 => (others => 237), 
171 => (others => 238), 
172 => (others => 239), 
173 => (others => 240), 
174 => (others => 241), 
175 => (others => 242), 
176 => (others => 243), 
177 => (others => 244), 
178 => (others => 245), 
179 => (others => 246), 
180 => (others => 247), 
181 => (others => 208), 
182 => (others => 209), 
183 => (others => 210), 
184 => (others => 238), 
185 => (others => 238), 
186 => (others => 239), 
187 => (others => 240), 
188 => (others => 241), 
189 => (others => 242), 
190 => (others => 242), 
191 => (others => 243), 
192 => (others => 243), 
193 => (others => 244), 
194 => (others => 245), 
195 => (others => 246), 
196 => (others => 247), 
197 => (others => 248), 
198 => (others => 251), 
199 => (others => 252), 
200 => (others => 253), 
201 => (others => 254), 
202 => (others => 255), 
203 => (others => 210), 
204 => (others => 211), 
205 => (others => 212), 
206 => (others => 213), 
207 => (others => 214), 
208 => (others => 215), 
209 => (others => 216), 
210 => (others => 217), 
211 => (others => 218), 
212 => (others => 219), 
213 => (others => 220), 
214 => (others => 221), 
215 => (others => 222), 
others => (others => 0)), others => (others => (others => 0))),
others => (others => (others => (others => 0))))
);
constant psi1_volt_LUT : voltage_LUT :=(
(15 => (7 => (0 => (others => 19), 
1 => (others => 19), 
2 => (others => 19), 
3 => (others => 20), 
4 => (others => 20), 
5 => (others => 20), 
6 => (others => 21), 
7 => (others => 21), 
8 => (others => 21), 
9 => (others => 21), 
10 => (others => 22), 
11 => (others => 22), 
12 => (others => 22), 
13 => (others => 22), 
14 => (others => 23), 
15 => (others => 23), 
16 => (others => 124), 
17 => (others => 124), 
18 => (others => 124), 
19 => (others => 125), 
20 => (others => 125), 
21 => (others => 125), 
22 => (others => 125), 
23 => (others => 125), 
24 => (others => 126), 
25 => (others => 126), 
26 => (others => 126), 
27 => (others => 126), 
28 => (others => 127), 
29 => (others => 127), 
30 => (others => 127), 
31 => (others => 127), 
32 => (others => 127), 
33 => (others => 127), 
34 => (others => 128), 
35 => (others => 145), 
36 => (others => 146), 
37 => (others => 146), 
38 => (others => 146), 
39 => (others => 146), 
40 => (others => 147), 
41 => (others => 147), 
42 => (others => 147), 
43 => (others => 147), 
44 => (others => 148), 
45 => (others => 143), 
46 => (others => 143), 
47 => (others => 143), 
48 => (others => 144), 
49 => (others => 144), 
50 => (others => 144), 
51 => (others => 145), 
52 => (others => 145), 
53 => (others => 145), 
54 => (others => 146), 
55 => (others => 146), 
56 => (others => 146), 
57 => (others => 147), 
58 => (others => 190), 
59 => (others => 190), 
60 => (others => 190), 
61 => (others => 190), 
62 => (others => 191), 
63 => (others => 191), 
64 => (others => 191), 
65 => (others => 192), 
66 => (others => 192), 
67 => (others => 192), 
68 => (others => 192), 
69 => (others => 193), 
70 => (others => 193), 
71 => (others => 193), 
72 => (others => 121), 
73 => (others => 121), 
74 => (others => 122), 
75 => (others => 122), 
76 => (others => 122), 
77 => (others => 123), 
78 => (others => 123), 
79 => (others => 157), 
80 => (others => 157), 
81 => (others => 158), 
82 => (others => 158), 
83 => (others => 158), 
84 => (others => 159), 
85 => (others => 159), 
86 => (others => 159), 
87 => (others => 160), 
88 => (others => 160), 
89 => (others => 160), 
90 => (others => 160), 
91 => (others => 161), 
92 => (others => 126), 
93 => (others => 126), 
94 => (others => 127), 
95 => (others => 127), 
96 => (others => 127), 
97 => (others => 127), 
98 => (others => 128), 
99 => (others => 128), 
100 => (others => 128), 
101 => (others => 129), 
102 => (others => 129), 
103 => (others => 129), 
104 => (others => 129), 
105 => (others => 130), 
106 => (others => 130), 
107 => (others => 145), 
108 => (others => 145), 
109 => (others => 145), 
110 => (others => 146), 
111 => (others => 146), 
112 => (others => 146), 
113 => (others => 147), 
114 => (others => 147), 
115 => (others => 208), 
116 => (others => 209), 
117 => (others => 209), 
118 => (others => 209), 
119 => (others => 209), 
120 => (others => 210), 
121 => (others => 210), 
122 => (others => 210), 
123 => (others => 211), 
124 => (others => 211), 
125 => (others => 211), 
126 => (others => 211), 
127 => (others => 212), 
128 => (others => 212), 
129 => (others => 212), 
130 => (others => 193), 
131 => (others => 193), 
132 => (others => 193), 
133 => (others => 194), 
134 => (others => 194), 
135 => (others => 194), 
136 => (others => 194), 
137 => (others => 195), 
138 => (others => 195), 
139 => (others => 195), 
140 => (others => 195), 
141 => (others => 196), 
142 => (others => 196), 
143 => (others => 196), 
144 => (others => 196), 
145 => (others => 196), 
146 => (others => 197), 
147 => (others => 175), 
148 => (others => 175), 
149 => (others => 175), 
150 => (others => 176), 
151 => (others => 126), 
152 => (others => 126), 
153 => (others => 126), 
154 => (others => 127), 
155 => (others => 127), 
156 => (others => 127), 
157 => (others => 128), 
158 => (others => 128), 
159 => (others => 128), 
160 => (others => 128), 
161 => (others => 129), 
162 => (others => 129), 
163 => (others => 129), 
164 => (others => 129), 
165 => (others => 130), 
166 => (others => 119), 
167 => (others => 119), 
168 => (others => 119), 
169 => (others => 41), 
170 => (others => 41), 
171 => (others => 41), 
172 => (others => 42), 
173 => (others => 42), 
174 => (others => 42), 
175 => (others => 43), 
176 => (others => 43), 
177 => (others => 43), 
178 => (others => 44), 
179 => (others => 44), 
180 => (others => 44), 
181 => (others => 143), 
182 => (others => 143), 
183 => (others => 143), 
184 => (others => 179), 
185 => (others => 180), 
186 => (others => 180), 
187 => (others => 180), 
188 => (others => 180), 
189 => (others => 181), 
190 => (others => 181), 
191 => (others => 181), 
192 => (others => 181), 
193 => (others => 181), 
194 => (others => 182), 
195 => (others => 182), 
196 => (others => 182), 
197 => (others => 183), 
198 => (others => 135), 
199 => (others => 135), 
200 => (others => 136), 
201 => (others => 136), 
202 => (others => 136), 
203 => (others => 210), 
204 => (others => 210), 
205 => (others => 210), 
206 => (others => 211), 
207 => (others => 211), 
208 => (others => 211), 
209 => (others => 212), 
210 => (others => 212), 
211 => (others => 212), 
212 => (others => 213), 
213 => (others => 213), 
214 => (others => 213), 
215 => (others => 213), 
others => (others => 0)), others => (others => (others => 0))),
others => (others => (others => (others => 0))))
);
constant psi2_volt_LUT : voltage_LUT :=(
(15 => (7 => (0 => (others => 140), 
1 => (others => 140), 
2 => (others => 141), 
3 => (others => 141), 
4 => (others => 141), 
5 => (others => 141), 
6 => (others => 141), 
7 => (others => 141), 
8 => (others => 141), 
9 => (others => 142), 
10 => (others => 142), 
11 => (others => 142), 
12 => (others => 142), 
13 => (others => 142), 
14 => (others => 142), 
15 => (others => 142), 
16 => (others => 201), 
17 => (others => 201), 
18 => (others => 201), 
19 => (others => 201), 
20 => (others => 201), 
21 => (others => 201), 
22 => (others => 201), 
23 => (others => 202), 
24 => (others => 202), 
25 => (others => 202), 
26 => (others => 202), 
27 => (others => 202), 
28 => (others => 202), 
29 => (others => 202), 
30 => (others => 202), 
31 => (others => 202), 
32 => (others => 202), 
33 => (others => 203), 
34 => (others => 203), 
35 => (others => 132), 
36 => (others => 132), 
37 => (others => 132), 
38 => (others => 132), 
39 => (others => 132), 
40 => (others => 132), 
41 => (others => 133), 
42 => (others => 133), 
43 => (others => 133), 
44 => (others => 133), 
45 => (others => 152), 
46 => (others => 152), 
47 => (others => 152), 
48 => (others => 153), 
49 => (others => 153), 
50 => (others => 153), 
51 => (others => 153), 
52 => (others => 153), 
53 => (others => 153), 
54 => (others => 154), 
55 => (others => 154), 
56 => (others => 154), 
57 => (others => 154), 
58 => (others => 172), 
59 => (others => 172), 
60 => (others => 172), 
61 => (others => 172), 
62 => (others => 172), 
63 => (others => 173), 
64 => (others => 173), 
65 => (others => 173), 
66 => (others => 173), 
67 => (others => 173), 
68 => (others => 173), 
69 => (others => 173), 
70 => (others => 174), 
71 => (others => 174), 
72 => (others => 95), 
73 => (others => 95), 
74 => (others => 95), 
75 => (others => 95), 
76 => (others => 95), 
77 => (others => 96), 
78 => (others => 96), 
79 => (others => 37), 
80 => (others => 37), 
81 => (others => 37), 
82 => (others => 37), 
83 => (others => 37), 
84 => (others => 37), 
85 => (others => 38), 
86 => (others => 38), 
87 => (others => 38), 
88 => (others => 38), 
89 => (others => 38), 
90 => (others => 38), 
91 => (others => 38), 
92 => (others => 127), 
93 => (others => 127), 
94 => (others => 127), 
95 => (others => 127), 
96 => (others => 128), 
97 => (others => 128), 
98 => (others => 128), 
99 => (others => 128), 
100 => (others => 128), 
101 => (others => 128), 
102 => (others => 128), 
103 => (others => 129), 
104 => (others => 129), 
105 => (others => 129), 
106 => (others => 129), 
107 => (others => 193), 
108 => (others => 193), 
109 => (others => 193), 
110 => (others => 194), 
111 => (others => 194), 
112 => (others => 194), 
113 => (others => 194), 
114 => (others => 194), 
115 => (others => 237), 
116 => (others => 237), 
117 => (others => 237), 
118 => (others => 237), 
119 => (others => 237), 
120 => (others => 238), 
121 => (others => 238), 
122 => (others => 238), 
123 => (others => 238), 
124 => (others => 238), 
125 => (others => 238), 
126 => (others => 239), 
127 => (others => 239), 
128 => (others => 239), 
129 => (others => 239), 
130 => (others => 161), 
131 => (others => 161), 
132 => (others => 161), 
133 => (others => 161), 
134 => (others => 161), 
135 => (others => 162), 
136 => (others => 162), 
137 => (others => 162), 
138 => (others => 162), 
139 => (others => 162), 
140 => (others => 162), 
141 => (others => 162), 
142 => (others => 162), 
143 => (others => 163), 
144 => (others => 163), 
145 => (others => 163), 
146 => (others => 163), 
147 => (others => 199), 
148 => (others => 199), 
149 => (others => 199), 
150 => (others => 199), 
151 => (others => 165), 
152 => (others => 165), 
153 => (others => 165), 
154 => (others => 165), 
155 => (others => 165), 
156 => (others => 165), 
157 => (others => 166), 
158 => (others => 166), 
159 => (others => 166), 
160 => (others => 166), 
161 => (others => 166), 
162 => (others => 166), 
163 => (others => 166), 
164 => (others => 166), 
165 => (others => 166), 
166 => (others => 194), 
167 => (others => 194), 
168 => (others => 194), 
169 => (others => 87), 
170 => (others => 87), 
171 => (others => 87), 
172 => (others => 87), 
173 => (others => 87), 
174 => (others => 87), 
175 => (others => 88), 
176 => (others => 88), 
177 => (others => 88), 
178 => (others => 88), 
179 => (others => 88), 
180 => (others => 88), 
181 => (others => 95), 
182 => (others => 95), 
183 => (others => 95), 
184 => (others => 14), 
185 => (others => 14), 
186 => (others => 14), 
187 => (others => 14), 
188 => (others => 14), 
189 => (others => 14), 
190 => (others => 15), 
191 => (others => 15), 
192 => (others => 15), 
193 => (others => 15), 
194 => (others => 15), 
195 => (others => 15), 
196 => (others => 15), 
197 => (others => 15), 
198 => (others => 20), 
199 => (others => 20), 
200 => (others => 20), 
201 => (others => 20), 
202 => (others => 20), 
203 => (others => 210), 
204 => (others => 210), 
205 => (others => 210), 
206 => (others => 210), 
207 => (others => 210), 
208 => (others => 210), 
209 => (others => 211), 
210 => (others => 211), 
211 => (others => 211), 
212 => (others => 211), 
213 => (others => 211), 
214 => (others => 211), 
215 => (others => 211), 
others => (others => 0)), others => (others => (others => 0))),
others => (others => (others => (others => 0))))
);
constant psi3_volt_LUT : voltage_LUT :=(
(15 => (7 => (0 => (others => 154), 
1 => (others => 155), 
2 => (others => 155), 
3 => (others => 155), 
4 => (others => 155), 
5 => (others => 155), 
6 => (others => 155), 
7 => (others => 155), 
8 => (others => 155), 
9 => (others => 155), 
10 => (others => 155), 
11 => (others => 155), 
12 => (others => 155), 
13 => (others => 155), 
14 => (others => 155), 
15 => (others => 155), 
16 => (others => 23), 
17 => (others => 23), 
18 => (others => 23), 
19 => (others => 23), 
20 => (others => 23), 
21 => (others => 23), 
22 => (others => 23), 
23 => (others => 23), 
24 => (others => 23), 
25 => (others => 23), 
26 => (others => 23), 
27 => (others => 23), 
28 => (others => 23), 
29 => (others => 23), 
30 => (others => 23), 
31 => (others => 23), 
32 => (others => 24), 
33 => (others => 24), 
34 => (others => 24), 
35 => (others => 92), 
36 => (others => 92), 
37 => (others => 92), 
38 => (others => 92), 
39 => (others => 92), 
40 => (others => 92), 
41 => (others => 92), 
42 => (others => 92), 
43 => (others => 92), 
44 => (others => 92), 
45 => (others => 249), 
46 => (others => 249), 
47 => (others => 249), 
48 => (others => 249), 
49 => (others => 249), 
50 => (others => 249), 
51 => (others => 249), 
52 => (others => 249), 
53 => (others => 249), 
54 => (others => 250), 
55 => (others => 250), 
56 => (others => 250), 
57 => (others => 250), 
58 => (others => 146), 
59 => (others => 146), 
60 => (others => 146), 
61 => (others => 146), 
62 => (others => 146), 
63 => (others => 146), 
64 => (others => 147), 
65 => (others => 147), 
66 => (others => 147), 
67 => (others => 147), 
68 => (others => 147), 
69 => (others => 147), 
70 => (others => 147), 
71 => (others => 147), 
72 => (others => 46), 
73 => (others => 46), 
74 => (others => 46), 
75 => (others => 46), 
76 => (others => 47), 
77 => (others => 47), 
78 => (others => 47), 
79 => (others => 140), 
80 => (others => 140), 
81 => (others => 141), 
82 => (others => 141), 
83 => (others => 141), 
84 => (others => 141), 
85 => (others => 141), 
86 => (others => 141), 
87 => (others => 141), 
88 => (others => 141), 
89 => (others => 141), 
90 => (others => 141), 
91 => (others => 141), 
92 => (others => 128), 
93 => (others => 128), 
94 => (others => 128), 
95 => (others => 128), 
96 => (others => 128), 
97 => (others => 128), 
98 => (others => 128), 
99 => (others => 128), 
100 => (others => 128), 
101 => (others => 128), 
102 => (others => 128), 
103 => (others => 128), 
104 => (others => 128), 
105 => (others => 128), 
106 => (others => 128), 
107 => (others => 77), 
108 => (others => 77), 
109 => (others => 77), 
110 => (others => 77), 
111 => (others => 77), 
112 => (others => 77), 
113 => (others => 77), 
114 => (others => 77), 
115 => (others => 65), 
116 => (others => 65), 
117 => (others => 65), 
118 => (others => 66), 
119 => (others => 66), 
120 => (others => 66), 
121 => (others => 66), 
122 => (others => 66), 
123 => (others => 66), 
124 => (others => 66), 
125 => (others => 66), 
126 => (others => 66), 
127 => (others => 66), 
128 => (others => 66), 
129 => (others => 66), 
130 => (others => 69), 
131 => (others => 69), 
132 => (others => 69), 
133 => (others => 69), 
134 => (others => 69), 
135 => (others => 69), 
136 => (others => 69), 
137 => (others => 69), 
138 => (others => 69), 
139 => (others => 69), 
140 => (others => 69), 
141 => (others => 69), 
142 => (others => 69), 
143 => (others => 69), 
144 => (others => 69), 
145 => (others => 70), 
146 => (others => 70), 
147 => (others => 119), 
148 => (others => 119), 
149 => (others => 119), 
150 => (others => 119), 
151 => (others => 202), 
152 => (others => 203), 
153 => (others => 203), 
154 => (others => 203), 
155 => (others => 203), 
156 => (others => 203), 
157 => (others => 203), 
158 => (others => 203), 
159 => (others => 203), 
160 => (others => 203), 
161 => (others => 203), 
162 => (others => 203), 
163 => (others => 203), 
164 => (others => 203), 
165 => (others => 203), 
166 => (others => 240), 
167 => (others => 240), 
168 => (others => 240), 
169 => (others => 151), 
170 => (others => 151), 
171 => (others => 151), 
172 => (others => 151), 
173 => (others => 151), 
174 => (others => 152), 
175 => (others => 152), 
176 => (others => 152), 
177 => (others => 152), 
178 => (others => 152), 
179 => (others => 152), 
180 => (others => 152), 
181 => (others => 234), 
182 => (others => 234), 
183 => (others => 234), 
184 => (others => 34), 
185 => (others => 34), 
186 => (others => 34), 
187 => (others => 34), 
188 => (others => 34), 
189 => (others => 34), 
190 => (others => 34), 
191 => (others => 34), 
192 => (others => 34), 
193 => (others => 34), 
194 => (others => 35), 
195 => (others => 35), 
196 => (others => 35), 
197 => (others => 35), 
198 => (others => 171), 
199 => (others => 171), 
200 => (others => 171), 
201 => (others => 171), 
202 => (others => 171), 
203 => (others => 210), 
204 => (others => 210), 
205 => (others => 210), 
206 => (others => 210), 
207 => (others => 210), 
208 => (others => 210), 
209 => (others => 210), 
210 => (others => 210), 
211 => (others => 210), 
212 => (others => 210), 
213 => (others => 210), 
214 => (others => 210), 
215 => (others => 210), 
others => (others => 0)), others => (others => (others => 0))),
others => (others => (others => (others => 0))))
);
constant psi4_volt_LUT : voltage_LUT :=(
(15 => (7 => (0 => (others => 56), 
1 => (others => 57), 
2 => (others => 57), 
3 => (others => 57), 
4 => (others => 57), 
5 => (others => 57), 
6 => (others => 57), 
7 => (others => 57), 
8 => (others => 57), 
9 => (others => 57), 
10 => (others => 57), 
11 => (others => 57), 
12 => (others => 57), 
13 => (others => 57), 
14 => (others => 57), 
15 => (others => 57), 
16 => (others => 23), 
17 => (others => 23), 
18 => (others => 23), 
19 => (others => 23), 
20 => (others => 23), 
21 => (others => 23), 
22 => (others => 23), 
23 => (others => 23), 
24 => (others => 23), 
25 => (others => 23), 
26 => (others => 23), 
27 => (others => 23), 
28 => (others => 23), 
29 => (others => 23), 
30 => (others => 23), 
31 => (others => 24), 
32 => (others => 24), 
33 => (others => 24), 
34 => (others => 24), 
35 => (others => 92), 
36 => (others => 93), 
37 => (others => 93), 
38 => (others => 93), 
39 => (others => 93), 
40 => (others => 93), 
41 => (others => 93), 
42 => (others => 93), 
43 => (others => 93), 
44 => (others => 93), 
45 => (others => 56), 
46 => (others => 56), 
47 => (others => 56), 
48 => (others => 56), 
49 => (others => 56), 
50 => (others => 56), 
51 => (others => 56), 
52 => (others => 56), 
53 => (others => 56), 
54 => (others => 56), 
55 => (others => 56), 
56 => (others => 56), 
57 => (others => 56), 
58 => (others => 44), 
59 => (others => 44), 
60 => (others => 45), 
61 => (others => 45), 
62 => (others => 45), 
63 => (others => 45), 
64 => (others => 45), 
65 => (others => 45), 
66 => (others => 45), 
67 => (others => 45), 
68 => (others => 45), 
69 => (others => 45), 
70 => (others => 45), 
71 => (others => 45), 
72 => (others => 16), 
73 => (others => 16), 
74 => (others => 16), 
75 => (others => 16), 
76 => (others => 16), 
77 => (others => 16), 
78 => (others => 16), 
79 => (others => 127), 
80 => (others => 127), 
81 => (others => 127), 
82 => (others => 127), 
83 => (others => 127), 
84 => (others => 127), 
85 => (others => 127), 
86 => (others => 127), 
87 => (others => 127), 
88 => (others => 127), 
89 => (others => 127), 
90 => (others => 127), 
91 => (others => 127), 
92 => (others => 128), 
93 => (others => 128), 
94 => (others => 128), 
95 => (others => 128), 
96 => (others => 128), 
97 => (others => 128), 
98 => (others => 128), 
99 => (others => 128), 
100 => (others => 128), 
101 => (others => 128), 
102 => (others => 128), 
103 => (others => 128), 
104 => (others => 128), 
105 => (others => 128), 
106 => (others => 128), 
107 => (others => 230), 
108 => (others => 230), 
109 => (others => 230), 
110 => (others => 230), 
111 => (others => 230), 
112 => (others => 231), 
113 => (others => 231), 
114 => (others => 231), 
115 => (others => 19), 
116 => (others => 19), 
117 => (others => 19), 
118 => (others => 19), 
119 => (others => 20), 
120 => (others => 20), 
121 => (others => 20), 
122 => (others => 20), 
123 => (others => 20), 
124 => (others => 20), 
125 => (others => 20), 
126 => (others => 20), 
127 => (others => 20), 
128 => (others => 20), 
129 => (others => 20), 
130 => (others => 219), 
131 => (others => 219), 
132 => (others => 219), 
133 => (others => 219), 
134 => (others => 219), 
135 => (others => 219), 
136 => (others => 219), 
137 => (others => 219), 
138 => (others => 219), 
139 => (others => 219), 
140 => (others => 219), 
141 => (others => 219), 
142 => (others => 219), 
143 => (others => 220), 
144 => (others => 220), 
145 => (others => 220), 
146 => (others => 220), 
147 => (others => 128), 
148 => (others => 128), 
149 => (others => 128), 
150 => (others => 128), 
151 => (others => 157), 
152 => (others => 157), 
153 => (others => 157), 
154 => (others => 157), 
155 => (others => 157), 
156 => (others => 157), 
157 => (others => 157), 
158 => (others => 157), 
159 => (others => 158), 
160 => (others => 158), 
161 => (others => 158), 
162 => (others => 158), 
163 => (others => 158), 
164 => (others => 158), 
165 => (others => 158), 
166 => (others => 121), 
167 => (others => 121), 
168 => (others => 121), 
169 => (others => 242), 
170 => (others => 242), 
171 => (others => 242), 
172 => (others => 242), 
173 => (others => 242), 
174 => (others => 242), 
175 => (others => 242), 
176 => (others => 242), 
177 => (others => 242), 
178 => (others => 242), 
179 => (others => 242), 
180 => (others => 242), 
181 => (others => 233), 
182 => (others => 233), 
183 => (others => 233), 
184 => (others => 17), 
185 => (others => 17), 
186 => (others => 17), 
187 => (others => 17), 
188 => (others => 17), 
189 => (others => 17), 
190 => (others => 17), 
191 => (others => 17), 
192 => (others => 18), 
193 => (others => 18), 
194 => (others => 18), 
195 => (others => 18), 
196 => (others => 18), 
197 => (others => 18), 
198 => (others => 59), 
199 => (others => 59), 
200 => (others => 59), 
201 => (others => 59), 
202 => (others => 59), 
203 => (others => 210), 
204 => (others => 210), 
205 => (others => 210), 
206 => (others => 210), 
207 => (others => 210), 
208 => (others => 210), 
209 => (others => 210), 
210 => (others => 210), 
211 => (others => 210), 
212 => (others => 210), 
213 => (others => 210), 
214 => (others => 210), 
215 => (others => 210), 
others => (others => 0)), others => (others => (others => 0))),
others => (others => (others => (others => 0))))
);
signal my_theta_LUT: theta_LUT :=(0 => -14124, 1 => -14020, 2 => -14005, 3 => -13882, 4 => -13789, 5 => -13697, 6 => -13574, 7 => -13482, 8 => -13390, 9 => -13375, 10 => -13252, 11 => -13160, 12 => -13068, 13 => -12977, 14 => -12946, 15 => -12854, 16 => -11564, 17 => -11473, 18 => -11381, 19 => -11351, 20 => -11260, 21 => -11168, 22 => -11077, 23 => -11062, 24 => -11032, 25 => -10940, 26 => -10849, 27 => -10758, 28 => -10728, 29 => -10637, 30 => -10546, 31 => -10542, 32 => -10443, 33 => -10428, 34 => -10398, 35 => -9912, 36 => -9878, 37 => -9788, 38 => -9697, 39 => -9606, 40 => -9576, 41 => -9470, 42 => -9379, 43 => -9288, 44 => -9258, 45 => -9254, 46 => -9164, 47 => -9073, 48 => -8937, 49 => -8846, 50 => -8756, 51 => -8635, 52 => -8544, 53 => -8454, 54 => -8311, 55 => -8220, 56 => -8130, 57 => -8009, 58 => -6640, 59 => -6550, 60 => -6456, 61 => -6366, 62 => -6246, 63 => -6141, 64 => -6043, 65 => -6013, 66 => -5923, 67 => -5833, 68 => -5743, 69 => -5623, 70 => -5519, 71 => -5429, 72 => -5320, 73 => -5230, 74 => -5110, 75 => -5020, 76 => -4923, 77 => -4878, 78 => -4788, 79 => -2467, 80 => -2377, 81 => -2250, 82 => -2161, 83 => -2071, 84 => -1952, 85 => -1847, 86 => -1758, 87 => -1638, 88 => -1549, 89 => -1459, 90 => -1370, 91 => -1340, 92 => -612, 93 => -523, 94 => -403, 95 => -314, 96 => -299, 97 => -209, 98 => -90, 99 => -1, 100 => 89, 101 => 208, 102 => 298, 103 => 313, 104 => 402, 105 => 522, 106 => 611, 107 => 671, 108 => 760, 109 => 850, 110 => 984, 111 => 1074, 112 => 1167, 113 => 1287, 114 => 1376, 115 => 1973, 116 => 2003, 117 => 2093, 118 => 2100, 119 => 2193, 120 => 2328, 121 => 2417, 122 => 2507, 123 => 2626, 124 => 2716, 125 => 2806, 126 => 2910, 127 => 2940, 128 => 3030, 129 => 3119, 130 => 3856, 131 => 3945, 132 => 4035, 133 => 4065, 134 => 4155, 135 => 4260, 136 => 4349, 137 => 4379, 138 => 4469, 139 => 4559, 140 => 4649, 141 => 4679, 142 => 4768, 143 => 4877, 144 => 4967, 145 => 4974, 146 => 5004, 147 => 5087, 148 => 5177, 149 => 5266, 150 => 5386, 151 => 5458, 152 => 5555, 153 => 5645, 154 => 5765, 155 => 5855, 156 => 5945, 157 => 6080, 158 => 6170, 159 => 6264, 160 => 6354, 161 => 6384, 162 => 6474, 163 => 6564, 164 => 6654, 165 => 6684, 166 => 6733, 167 => 6823, 168 => 6913, 169 => 7075, 170 => 7165, 171 => 7255, 172 => 7376, 173 => 7466, 174 => 7564, 175 => 7699, 176 => 7790, 177 => 7880, 178 => 8001, 179 => 8091, 180 => 8181, 181 => 8328, 182 => 8419, 183 => 8509, 184 => 8585, 185 => 8615, 186 => 8706, 187 => 8796, 188 => 8887, 189 => 9008, 190 => 9023, 191 => 9113, 192 => 9117, 193 => 9208, 194 => 9336, 195 => 9427, 196 => 9518, 197 => 9639, 198 => 9718, 199 => 9809, 200 => 9930, 201 => 10021, 202 => 10112, 203 => 12017, 204 => 12108, 205 => 12200, 206 => 12322, 207 => 12413, 208 => 12505, 209 => 12643, 210 => 12735, 211 => 12826, 212 => 12949, 213 => 13041, 214 => 13133, 215 => 13225, others=>0);
begin    
    updater : process(clk) begin
        if rising_edge(clk) then
            necessary_voltage_psi0 <= psi0_volt_LUT(requested_row,requested_col,requested_theta,requested_phi);
            necessary_voltage_psi1 <= psi1_volt_LUT(requested_row,requested_col,requested_theta,requested_phi);
            necessary_voltage_psi2 <= psi2_volt_LUT(requested_row,requested_col,requested_theta,requested_phi);
            necessary_voltage_psi3 <= psi3_volt_LUT(requested_row,requested_col,requested_theta,requested_phi);
            necessary_voltage_psi4 <= psi4_volt_LUT(requested_row,requested_col,requested_theta,requested_phi);
            returned_theta_ang <= my_theta_LUT(requested_theta);
        end if;
    end process;

end Behavioral;