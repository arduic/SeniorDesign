package fft_len is
constant LOG2_FFT_LEN: integer := 10;
constant FFT_LEN: integer := 1024;
constant ICPX_WIDTH: integer := 16;
constant INPUT_FILE: string := "C:\Users\lc599.DREXEL\SeniorDesign\FFT\scripts\data_in.txt";
constant OUTPUT_FILE: string := "C:\Users\lc599.DREXEL\SeniorDesign\FFT\scripts\data_out.txt";
end fft_len;
